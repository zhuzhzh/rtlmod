module udp_dff();
reg a;
endmodule
