module udp_sedfft();
reg a;
endmodule
